module decoder_4_to_16(
	input wire [3:0] a,
	output reg [15:0] b
);
always @(*)
begin
    case (a)
		 4'b0000 : b <= 16'b0000000000000001;
		 4'b0001 : b <= 16'b0000000000000010;
		 4'b0010 : b <= 16'b0000000000000100;
		 4'b0011 : b <= 16'b0000000000001000;
		 4'b0100 : b <= 16'b0000000000010000;
		 4'b0101 : b <= 16'b0000000000100000;
		 4'b0110 : b <= 16'b0000000001000000;
		 4'b0111 : b <= 16'b0000000010000000;
		 4'b1000 : b <= 16'b0000000100000000;
		 4'b1001 : b <= 16'b0000001000000000;
		 4'b1010 : b <= 16'b0000010000000000;
		 4'b1011 : b <= 16'b0000100000000000;
		 4'b1100 : b <= 16'b0001000000000000;
		 4'b1101 : b <= 16'b0010000000000000;
		 4'b1110 : b <= 16'b0100000000000000;
		 4'b1111 : b <= 16'b1000000000000000;
		 default : b <= 16'b0000000000000000;
	 endcase
end
endmodule
	 
	 
	 